// D4
// test send in
/*
   author: jc21g13
   last revision: 01 Mar' 15
*/

module test_data(output logic[7:0] data);

assign data = 8'b01001001;

endmodule 